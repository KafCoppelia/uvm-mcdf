`ifndef TRANSACTION_PKG_SV
`define TRANSACTION_PKG_SV

`include "transaction_channel.sv"
`include "transaction_bus.sv"
`include "transaction_formater.sv"

`endif

