`ifndef AGENT_PKG_SV
`define AGENT_PKG_SV

`include "agent_bus.sv"
`include "agent_channel.sv"
`include "agent_formater.sv"
`include "agent_pkg.sv"

`endif

