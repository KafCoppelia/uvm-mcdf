`ifndef MONITOR_PKG_SV
`define MONITOR_PKG_SV

`include "monitor_bus.sv"
`include "monitor_channel.sv"
`include "monitor_formater.sv"

`endif

