`ifndef REGISTER_PKG_SV
`define REGISTER_PKG_SV

`include "adapter.sv"
`include "reg_model.sv"

`endif

